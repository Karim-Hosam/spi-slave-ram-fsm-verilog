module SPI_Slave_with_Ram(
    port_list
);
    
endmodule