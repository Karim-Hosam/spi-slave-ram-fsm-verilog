module SPI_Slave(
    port_list
);
    
endmodule