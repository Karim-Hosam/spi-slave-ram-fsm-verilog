module Counter(
    input clk;
    input reset,
    input enable,
);
    
endmodule