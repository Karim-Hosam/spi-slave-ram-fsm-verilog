module Single_Port_Sync_RAM(
    port_list
);
    
endmodule