module SPI_Slave_with_Ram_tb(
    port_list
);
    
endmodule